module title(
    input  wire       clk,
    input  wire [7:0] ascii,
    input  wire [3:0] row,
    output reg  [7:0] pixels
);

    reg [7:0] font[0:128*8-1];

    initial begin
        //B
        font["B"*8+0] = 8'b11111100;
        font["B"*8+1] = 8'b11000110;
        font["B"*8+2] = 8'b11000110;
        font["B"*8+3] = 8'b11111100;
        font["B"*8+4] = 8'b11000110;
        font["B"*8+5] = 8'b11000110;
        font["B"*8+6] = 8'b11111100;
        font["B"*8+7] = 8'b00000000;

        //R
        font["R"*8+0] = 8'b11111100;
        font["R"*8+1] = 8'b11000110;
        font["R"*8+2] = 8'b11000110;
        font["R"*8+3] = 8'b11111100;
        font["R"*8+4] = 8'b11100000;
        font["R"*8+5] = 8'b11011000;
        font["R"*8+6] = 8'b11001100;
        font["R"*8+7] = 8'b00000000;

        //E
        font["E"*8+0] = 8'b11111110;
        font["E"*8+1] = 8'b11000000;
        font["E"*8+2] = 8'b11000000;
        font["E"*8+3] = 8'b11111100;
        font["E"*8+4] = 8'b11000000;
        font["E"*8+5] = 8'b11000000;
        font["E"*8+6] = 8'b11111110;
        font["E"*8+7] = 8'b00000000;

        //A
        font["A"*8+0] = 8'b01111100;
        font["A"*8+1] = 8'b11000110;
        font["A"*8+2] = 8'b11000110;
        font["A"*8+3] = 8'b11111110;
        font["A"*8+4] = 8'b11000110;
        font["A"*8+5] = 8'b11000110;
        font["A"*8+6] = 8'b11000110;
        font["A"*8+7] = 8'b00000000;

        //K
        font["K"*8+0] = 8'b11000110;
        font["K"*8+1] = 8'b11001100;
        font["K"*8+2] = 8'b11011000;
        font["K"*8+3] = 8'b11110000;
        font["K"*8+4] = 8'b11110000;
        font["K"*8+5] = 8'b11011000;
        font["K"*8+6] = 8'b11001100;
        font["K"*8+7] = 8'b00000000;

        //O
        font["O"*8+0] = 8'b01111100;
        font["O"*8+1] = 8'b11000110;
        font["O"*8+2] = 8'b11000110;
        font["O"*8+3] = 8'b11000110;
        font["O"*8+4] = 8'b11000110;
        font["O"*8+5] = 8'b11000110;
        font["O"*8+6] = 8'b01111100;
        font["O"*8+7] = 8'b00000000;

        //U
        font["U"*8+0] = 8'b11000110;
        font["U"*8+1] = 8'b11000110;
        font["U"*8+2] = 8'b11000110;
        font["U"*8+3] = 8'b11000110;
        font["U"*8+4] = 8'b11000110;
        font["U"*8+5] = 8'b11000110;
        font["U"*8+6] = 8'b01111100;
        font["U"*8+7] = 8'b00000000;

        //T
        font["T"*8+0] = 8'b11111110;
        font["T"*8+1] = 8'b00110000;
        font["T"*8+2] = 8'b00110000;
        font["T"*8+3] = 8'b00110000;
        font["T"*8+4] = 8'b00110000;
        font["T"*8+5] = 8'b00110000;
        font["T"*8+6] = 8'b00110000;
        font["T"*8+7] = 8'b00000000;

        //S
        font["S"*8+0] = 8'b01111110;
        font["S"*8+1] = 8'b11000000;
        font["S"*8+2] = 8'b11000000;
        font["S"*8+3] = 8'b01111100;
        font["S"*8+4] = 8'b00000110;
        font["S"*8+5] = 8'b00000110;
        font["S"*8+6] = 8'b11111100;
        font["S"*8+7] = 8'b00000000;

        //L
        font["L"*8+0] = 8'b11000000;
        font["L"*8+1] = 8'b11000000;
        font["L"*8+2] = 8'b11000000;
        font["L"*8+3] = 8'b11000000;
        font["L"*8+4] = 8'b11000000;
        font["L"*8+5] = 8'b11000000;
        font["L"*8+6] = 8'b11111110;
        font["L"*8+7] = 8'b00000000;

        //F
        font["F"*8+0] = 8'b11111110;
        font["F"*8+1] = 8'b11000000;
        font["F"*8+2] = 8'b11000000;
        font["F"*8+3] = 8'b11111100;
        font["F"*8+4] = 8'b11000000;
        font["F"*8+5] = 8'b11000000;
        font["F"*8+6] = 8'b11000000;
        font["F"*8+7] = 8'b00000000;

        //G
        font["G"*8+0] = 8'b01111100;
        font["G"*8+1] = 8'b11000110;
        font["G"*8+2] = 8'b11000000;
        font["G"*8+3] = 8'b11000000;
        font["G"*8+4] = 8'b11001110;
        font["G"*8+5] = 8'b11000110;
        font["G"*8+6] = 8'b01111100;
        font["G"*8+7] = 8'b00000000;

        //H
        font["H"*8+0] = 8'b11000110;
        font["H"*8+1] = 8'b11000110;
        font["H"*8+2] = 8'b11000110;
        font["H"*8+3] = 8'b11111110;
        font["H"*8+4] = 8'b11000110;
        font["H"*8+5] = 8'b11000110;
        font["H"*8+6] = 8'b11000110;
        font["H"*8+7] = 8'b00000000;

        //P
        font["P"*8+0] = 8'b11111100;
        font["P"*8+1] = 8'b11000110;
        font["P"*8+2] = 8'b11000110;
        font["P"*8+3] = 8'b11111100;
        font["P"*8+4] = 8'b11000000;
        font["P"*8+5] = 8'b11000000;
        font["P"*8+6] = 8'b11000000;
        font["P"*8+7] = 8'b00000000;

        //Y
        font["Y"*8+0] = 8'b11000110;
        font["Y"*8+1] = 8'b11000110;
        font["Y"*8+2] = 8'b01101100;
        font["Y"*8+3] = 8'b00111000;
        font["Y"*8+4] = 8'b00111000;
        font["Y"*8+5] = 8'b00111000;
        font["Y"*8+6] = 8'b00111000;
        font["Y"*8+7] = 8'b00000000;
		  
		  //W
		  font["W"*8+0] = 8'b11000110;
		  font["W"*8+1] = 8'b11000110;
		  font["W"*8+2] = 8'b11000110;
		  font["W"*8+3] = 8'b11010110;
		  font["W"*8+4] = 8'b11111110;
		  font["W"*8+5] = 8'b11101110;
		  font["W"*8+6] = 8'b11000110;
		  font["W"*8+7] = 8'b00000000;

			//I
		  font["I"*8+0] = 8'b11111110;
		  font["I"*8+1] = 8'b00110000;
		  font["I"*8+2] = 8'b00110000;
		  font["I"*8+3] = 8'b00110000;
		  font["I"*8+4] = 8'b00110000;
		  font["I"*8+5] = 8'b00110000;
		  font["I"*8+6] = 8'b11111110;
		  font["I"*8+7] = 8'b00000000;

        //1
        font["1"*8+0] = 8'b00011000;
        font["1"*8+1] = 8'b00111000;
        font["1"*8+2] = 8'b00011000;
        font["1"*8+3] = 8'b00011000;
        font["1"*8+4] = 8'b00011000;
        font["1"*8+5] = 8'b00011000;
        font["1"*8+6] = 8'b01111110;
        font["1"*8+7] = 8'b00000000;
		  
		  // 2
		  font["2"*8+0] = 8'b00111100;
		  font["2"*8+1] = 8'b01111110;
		  font["2"*8+2] = 8'b11000110;
		  font["2"*8+3] = 8'b00001100;
		  font["2"*8+4] = 8'b00011000;
		  font["2"*8+5] = 8'b00110000;
		  font["2"*8+6] = 8'b01111110;
		  font["2"*8+7] = 8'b00000000;


        //3
        font["3"*8+0] = 8'b01111100;
        font["3"*8+1] = 8'b11000110;
        font["3"*8+2] = 8'b00000110;
        font["3"*8+3] = 8'b00111100;
        font["3"*8+4] = 8'b00000110;
        font["3"*8+5] = 8'b11000110;
        font["3"*8+6] = 8'b01111100;
        font["3"*8+7] = 8'b00000000;

        //4
        font["4"*8+0] = 8'b00011100;
        font["4"*8+1] = 8'b00111100;
        font["4"*8+2] = 8'b01101100;
        font["4"*8+3] = 8'b11001100;
        font["4"*8+4] = 8'b11111110;
        font["4"*8+5] = 8'b00001100;
        font["4"*8+6] = 8'b00001100;
        font["4"*8+7] = 8'b00000000;

        //:
        font[":"*8+0] = 8'b00000000;
        font[":"*8+1] = 8'b00011000;
        font[":"*8+2] = 8'b00011000;
        font[":"*8+3] = 8'b00000000;
        font[":"*8+4] = 8'b00011000;
        font[":"*8+5] = 8'b00011000;
        font[":"*8+6] = 8'b00000000;
        font[":"*8+7] = 8'b00000000;

        //space
        font[" "*8+0] = 8'b00000000;
        font[" "*8+1] = 8'b00000000;
        font[" "*8+2] = 8'b00000000;
        font[" "*8+3] = 8'b00000000;
        font[" "*8+4] = 8'b00000000;
        font[" "*8+5] = 8'b00000000;
        font[" "*8+6] = 8'b00000000;
        font[" "*8+7] = 8'b00000000;
		  
		  //:)
		  font[")"*8+0] = 8'b00111100;
		  font[")"*8+1] = 8'b01000010;
		  font[")"*8+2] = 8'b10100101;
		  font[")"*8+3] = 8'b10000001;
		  font[")"*8+4] = 8'b10100101;
		  font[")"*8+5] = 8'b10011001;
		  font[")"*8+6] = 8'b01000010;
	     font[")"*8+7] = 8'b00111100;
			
		  //N
		  font["N"*8+0] = 8'b11000010;
		  font["N"*8+1] = 8'b11100010;
		  font["N"*8+2] = 8'b11010010;
		  font["N"*8+3] = 8'b11001010;
		  font["N"*8+4] = 8'b11000110;
		  font["N"*8+5] = 8'b11000010;
		  font["N"*8+6] = 8'b11000010;
		  font["N"*8+7] = 8'b00000000;

		  //right arrow
		  font["*"*8+0] = 8'b00011000; 
		  font["*"*8+1] = 8'b00001100;
		  font["*"*8+2] = 8'b00000110;
		  font["*"*8+3] = 8'b11111111;
		  font["*"*8+4] = 8'b11111111;
		  font["*"*8+5] = 8'b00000110;
		  font["*"*8+6] = 8'b00001100;
		  font["*"*8+7] = 8'b00011000;

		  //?
		  font["?"*8+0] = 8'b00111100;
		  font["?"*8+1] = 8'b01000010;
		  font["?"*8+2] = 8'b00000100;
		  font["?"*8+3] = 8'b00001000;
		  font["?"*8+4] = 8'b00010000;
		  font["?"*8+5] = 8'b00000000;
		  font["?"*8+6] = 8'b00010000;
		  font["?"*8+7] = 8'b00000000;


    end

    always @(posedge clk)
        pixels <= font[ascii*8 + row];

endmodule
